module dac_out(
    input wire pwm_clk,
    input wire rst_n,
    input wire [11:0] din,
    output wire pwm_out
);

    获取完整代码，搜索闲鱼会员名：tb49263172

endmodule