module i2s_top(
    input clk,
    input rst_n,
    output reg [23:0] ldata,
    output reg [23:0] rdata,
    output ready,

    output mic_sck,
    output mic_ws,
    input mic_sd
);

    获取完整代码，搜索闲鱼会员名：tb49263172

endmodule
