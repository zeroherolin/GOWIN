`timescale 1ns/1ps

module sim_top();

    获取完整代码，搜索闲鱼会员名：tb49263172

endmodule