library verilog;
use verilog.vl_types.all;
entity sim_top is
end sim_top;
