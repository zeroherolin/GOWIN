module top(
    input clk27M,
    input rst_n,

    output mic_sck,
    output mic_ws,
    input mic_sd,

    output mic_out
);

    获取完整代码，搜索闲鱼会员名：tb49263172

endmodule